// Verilog code for XNOR Gate
module xnorGate (a, b, out);

input a, b;
output out;
assign out = ~(a ^ b);

endmodule
