// Verilog code for NOT Gate
module notGate (a, out);

input a;
output out;
assign out = ~a;

endmodule
